module d_flipflop(
    input clk,
    input rst,
    input d,
    output reg q
);


initial begin q <= 1'b0;   end 
always @(posedge clk ) begin
    if (rst)
        q <= 1'b0;
    else
        q <= d;
end

endmodule
